module madd #(
    parameters
) (
    ports
);
    
endmodule